@00000000
73 00 10 00 73 00 10 00 73 00 10 00 73 00 10 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
