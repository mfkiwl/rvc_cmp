@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 81 00 00 93 81 00 00 13 82 00 00
93 82 00 00 13 83 00 00 93 83 00 00 13 84 00 00
93 84 00 00 13 85 00 00 93 85 00 00 13 86 00 00
93 86 00 00 13 87 00 00 93 87 00 00 13 88 00 00
93 88 00 00 13 89 00 00 93 89 00 00 13 8A 00 00
93 8A 00 00 13 8B 00 00 93 8B 00 00 13 8C 00 00
93 8C 00 00 13 8D 00 00 93 8D 00 00 13 8E 00 00
93 8E 00 00 13 8F 00 00 93 8F 00 00 93 00 10 00
13 01 20 00 93 01 30 00 13 05 00 40 23 20 15 00
23 22 25 00 23 24 35 00 03 22 05 00 83 22 45 00
03 23 85 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 73 00 10 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00
