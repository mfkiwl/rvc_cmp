@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 81 00 00 93 81 00 00 13 82 00 00
93 82 00 00 13 83 00 00 93 83 00 00 13 84 00 00
93 84 00 00 13 85 00 00 93 85 00 00 13 86 00 00
93 86 00 00 13 87 00 00 93 87 00 00 13 88 00 00
93 88 00 00 13 89 00 00 93 89 00 00 13 8A 00 00
93 8A 00 00 13 8B 00 00 93 8B 00 00 13 8C 00 00
93 8C 00 00 13 8D 00 00 93 8D 00 00 13 8E 00 00
93 8E 00 00 13 8F 00 00 93 8F 00 00 93 00 10 00
13 01 20 00 93 01 30 00 13 02 40 00 93 02 50 00
13 03 60 00 93 03 70 00 13 04 80 00 B3 24 11 00
33 B5 20 00 B3 55 12 00 33 F6 71 00 B3 16 11 00
33 87 40 00 B3 C7 51 00 33 E8 60 00 93 0F 00 40
23 20 15 00 23 22 25 00 23 24 35 00 23 26 45 00
23 28 55 00 23 2A 65 00 23 2C 75 00 23 2E 85 00
23 20 95 02 23 22 A5 02 23 24 B5 02 23 26 C5 02
23 28 D5 02 23 2A E5 02 23 2C F5 02 23 2E 05 03
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
73 00 10 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00
